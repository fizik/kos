component mosquitto.Setcommand

endpoints {
    setcommand : mosquitto.Setcommand
}